`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"

class environment;
  
  //generator and driver instance
  generator gen;
  driver    driv;
  monitor   	mon;
  scoreboard	scb;
  
  //mailbox handle's
  mailbox gen2driv;
  mailbox mon2scb;
  
  //virtual interface
  virtual ALU_intf vif;
  
  //constructor
  function new(virtual ALU_intf vif);
    //get the interface from test
    this.vif = vif;
    
    //creating the mailbox (Same handle will be shared across generator and driver)
    gen2driv = new();
    mon2scb  = new();
    
    //creating generator and driver
    gen  = new(gen2driv);
    driv = new(vif,gen2driv);
    mon  = new(vif,mon2scb);
    scb  = new(mon2scb);
  endfunction
  

  task pre_test();
    driv.reset();
  endtask
  
  task test();
    fork 
      gen.main();
      driv.main();
      mon.main();
      scb.main();
    join_any
  endtask
  
  task post_test();
    wait(gen.ended.triggered);
    
    wait(gen.count == driv.no_transactions);
    transaction_check: assert(gen.count == driv.no_transactions)
      $display("No of generation is equal to no of transaction in driver");
    else
      $error("No of generation is not equal to no of transaction in driver");
    
    wait(gen.count == scb.no_transactions);
    transaction_check2: assert(gen.count == scb.no_transactions)
      $display("No of generation is equal to no of transaction in scoreboard");
    else
      $error("No of generation is not equal to no of transaction in driver");
    
  endtask  
  
  //run task
  task run;
    pre_test();
    test();
    post_test();
    $finish;
  endtask
  
endclass
  
